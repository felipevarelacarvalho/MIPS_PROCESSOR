--MEM/WB