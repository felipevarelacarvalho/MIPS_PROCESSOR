--ID/EX