--EX/MEM