--IF/ID